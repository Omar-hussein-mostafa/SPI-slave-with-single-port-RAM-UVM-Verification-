module SLAVE (MOSI,MISO,SS_n,clk,rst_n,rx_data,rx_valid,tx_data,tx_valid);

localparam IDLE      = 3'b000;
localparam WRITE     = 3'b010;
localparam CHK_CMD   = 3'b001;
localparam READ_ADD  = 3'b011;
localparam READ_DATA = 3'b100;

input            MOSI, clk, rst_n, SS_n, tx_valid;
input      [7:0] tx_data;
output reg [9:0] rx_data;
output reg       rx_valid, MISO;

reg [3:0] counter;
reg       received_address;

reg [2:0] cs, ns;

always @(posedge clk) begin
    if (~rst_n) begin
        cs <= IDLE;
    end
    else begin
        cs <= ns;
    end
end

always @(*) begin
    case (cs)
        IDLE : begin
            if (SS_n)
                ns = IDLE;
            else
                ns = CHK_CMD;
        end
        CHK_CMD : begin
            if (SS_n)
                ns = IDLE;
            else begin
                if (~MOSI)
                    ns = WRITE;
                else begin
                    if (!received_address)          //Design Error : should check for not finishing Read_add 
                        ns = READ_ADD; 
                    else
                        ns = READ_DATA;
                end
            end
        end
        WRITE : begin
            if (SS_n)
                ns = IDLE;
            else
                ns = WRITE;
        end
        READ_ADD : begin
            if (SS_n)
                ns = IDLE;
            else
                ns = READ_ADD;
        end
        READ_DATA : begin
            if (SS_n)
                ns = IDLE;
            else
                ns = READ_DATA;
        end
    endcase
end

always @(posedge clk) begin
    if (~rst_n) begin 
        rx_data <= 0;
        rx_valid <= 0;
        received_address <= 0;
        MISO <= 0;
    end
    else begin
        case (cs)
            IDLE : begin
                rx_valid <= 0;
                MISO     <= 0;      //Design Error: MISO must be reseted 
                rx_data  <= 0;      //Design Error: should reset the rx_data

            end
            CHK_CMD : begin
                counter <= 10;      
            end
            WRITE : begin
                if (counter > 0) begin
                    rx_data[counter-1] <= MOSI;
                    counter <= counter - 1;
                end
                else begin
                    rx_valid <= 1;
                end
            end
            READ_ADD : begin
                if (counter > 0) begin
                    rx_data[counter-1] <= MOSI;
                    counter <= counter - 1;
                end
                else begin
                    rx_valid <= 1;
                    received_address <= 1;
                end
            end
            READ_DATA : begin
                if (tx_valid) begin
                    rx_valid <= 0;
                    if (counter > 0) begin
                        MISO <= tx_data[counter-1];
                        counter <= counter - 1;
                    end
                    else begin
                        MISO<=0;
                        received_address <= 0;
                    end
                end
                else begin
                    MISO<=0;
                    if (counter > 0) begin
                        rx_data[counter-1] <= MOSI;
                        counter <= counter - 1;
                    end
                    else begin
                        rx_valid <= 1;
                        counter <= 9;     //Design Error: the counter should be reloaded to 9 as the slave would wait one cycle for the tx_valid
                    end
                end
            end
        endcase
    end
end

`ifdef SIM
assert property(@(posedge clk) disable iff(!rst_n) (!SS_n && cs==IDLE) |-> ##1 cs==CHK_CMD);
assert property(@(posedge clk) disable iff(!rst_n) cs==CHK_CMD  |-> ##1 (cs==WRITE || cs==READ_ADD || cs==READ_DATA));
assert property(@(posedge clk) disable iff(!rst_n) cs==READ_ADD && $past(cs)==CHK_CMD |-> ##12 cs==IDLE);
assert property(@(posedge clk) disable iff(!rst_n) cs==READ_DATA && $past(cs)==CHK_CMD |-> ##22 cs==IDLE);
cover  property(@(posedge clk) disable iff(!rst_n) (!SS_n && cs==IDLE) |-> ##1 cs==CHK_CMD);
cover  property(@(posedge clk) disable iff(!rst_n) cs==CHK_CMD  |-> ##1 (cs==WRITE || cs==READ_ADD || cs==READ_DATA));
cover  property(@(posedge clk) disable iff(!rst_n) cs==READ_ADD && $past(cs)==CHK_CMD |-> ##12 cs==IDLE);
cover  property(@(posedge clk) disable iff(!rst_n) cs==READ_DATA && $past(cs)==CHK_CMD |-> ##22 cs==IDLE);
`endif 

endmodule