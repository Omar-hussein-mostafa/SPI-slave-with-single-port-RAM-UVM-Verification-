interface wrapper_if(clk);
    input clk;
    logic SS_n,rst_n,MOSI,MISO,MISO_exp;
endinterface