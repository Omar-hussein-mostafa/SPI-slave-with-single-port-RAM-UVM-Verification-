module RAM (din,clk,rst_n,rx_valid,dout,tx_valid);

input      [9:0] din;
input            clk, rst_n, rx_valid;

output reg [7:0] dout;
output reg       tx_valid;

reg [7:0] MEM [255:0];

reg [7:0] Rd_Addr, Wr_Addr;

always @(posedge clk) begin
    if (~rst_n) begin
        dout <= 0;
        tx_valid <= 0;
        Rd_Addr <= 0;
        Wr_Addr <= 0;
    end
    else  begin             //Design Error: missing begin and end
        if (rx_valid) begin
            case (din[9:8])
                2'b00 : Wr_Addr <= din[7:0];
                2'b01 : MEM[Wr_Addr] <= din[7:0];
                2'b10 : Rd_Addr <= din[7:0];
                2'b11 : dout <= MEM[Rd_Addr];           //Design Error : should be of Rd_addr
                default : dout <= 0;
            endcase
        end
        if(din[9] && din[8] && rx_valid) begin
            tx_valid<=1;
        end
        else if ((!din[9] || !din[8]) && rx_valid) begin
            tx_valid<=0;
        end
        //tx_valid <= (din[9] && din[8] && rx_valid)? 1'b1: 1'b0;
    end
end

endmodule